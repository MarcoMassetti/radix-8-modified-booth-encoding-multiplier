//Adder Unit

module au (
    input [25:0] G [8:0],	//Partial products
    input N [7:0], 			//Signs from both encoders
    output [47:0] Z);		//Sum


	//******FIRST LAYER******
	
    wire [31:21] s0_0;	//Sum outputs of the compressors (inputs of the next layer)
    wire [32:22] c0_0;	//Carry out of the compressors (inputs of the next layer)

    HA c0_21 (.A(G[0][21]), .B(G[1][21-3]), .S(s0_0[21]), .Co(c0_0[21+1]));
    HA c0_22 (.A(G[0][22]), .B(G[1][22-3]), .S(s0_0[22]), .Co(c0_0[22+1]));
    HA c0_23 (.A(G[0][23]), .B(G[1][23-3]), .S(s0_0[23]), .Co(c0_0[23+1]));
    FA c0_24(.A(G[0][24]), .B(G[1][24-3]), .Ci(G[2][24-6]),  .S(s0_0[24]), .Co(c0_0[24+1]));
    FA c0_25(.A(G[0][25]), .B(G[1][25-3]), .Ci(G[2][25-6]),  .S(s0_0[25]), .Co(c0_0[25+1]));
    FA c0_26(.A(N[0]), .B(G[1][26-3]), .Ci(G[2][26-6]),  .S(s0_0[26]), .Co(c0_0[26+1]));
    FA c0_27(.A(N[0]), .B(G[1][27-3]), .Ci(G[2][27-6]),  .S(s0_0[27]), .Co(c0_0[27+1]));
    FA c0_28(.A(N[0]), .B(G[1][28-3]), .Ci(G[2][28-6]),  .S(s0_0[28]), .Co(c0_0[28+1]));
    FA c0_29(.A(~N[0]), .B(~N[1]), .Ci(G[2][29-6]),  .S(s0_0[29]), .Co(c0_0[29+1]));
    HA c0_30 (.A(1'b1), .B(G[2][30-6]), .S(s0_0[30]), .Co(c0_0[30+1]));
    HA c0_31 (.A(1'b1), .B(G[2][31-6]), .S(s0_0[31]), .Co(c0_0[31+1]));


	//******FIRST ROW OF COMPRESSORS IN THE SECOND LAYER******

    wire [40:12] s1_0;	//Sum outputs of the compressors (inputs of the next layer)
    wire [41:13] c1_0;	//Carry out of the compressors (inputs of the next layer)
    wire [38:16] t1;	//Intermediate T between compressors of te same layer

    HA c1_12 (.A(G[0][12]), .B(G[1][12-3]), .S(s1_0[12]), .Co(c1_0[12+1]));
    HA c1_13 (.A(G[0][13]), .B(G[1][13-3]), .S(s1_0[13]), .Co(c1_0[13+1]));
    HA c1_14 (.A(G[0][14]), .B(G[1][14-3]), .S(s1_0[14]), .Co(c1_0[14+1]));
    Comp_4to2 c1_15(.X1(G[0][15]), .X2(G[1][15-3]), .X3(G[2][15-6]), .Ti(G[3][15-9]),  .S(s1_0[15]), .C(c1_0[15+1]), .To(t1[15+1]));
    Comp_4to2 c1_16(.X1(G[0][16]), .X2(G[1][16-3]), .X3(G[2][16-6]), .Ti(t1[15+1]),  .S(s1_0[16]), .C(c1_0[16+1]), .To(t1[16+1]));
    Comp_4to2 c1_17(.X1(G[0][17]), .X2(G[1][17-3]), .X3(G[2][17-6]), .Ti(t1[16+1]),  .S(s1_0[17]), .C(c1_0[17+1]), .To(t1[17+1]));
    Comp_5to3 c1_18(.X1(G[0][18]), .X2(G[1][18-3]), .X3(G[2][18-6]), .X4(G[3][18-9]), .Ti(t1[17+1]),  .S(s1_0[18]), .C(c1_0[18+1]), .To(t1[18+1]));
    Comp_5to3 c1_19(.X1(G[0][19]), .X2(G[1][19-3]), .X3(G[2][19-6]), .X4(G[3][19-9]), .Ti(t1[18+1]),  .S(s1_0[19]), .C(c1_0[19+1]), .To(t1[19+1]));
    Comp_5to3 c1_20(.X1(G[0][20]), .X2(G[1][20-3]), .X3(G[2][20-6]), .X4(G[3][20-9]), .Ti(t1[19+1]),  .S(s1_0[20]), .C(c1_0[20+1]), .To(t1[20+1]));
    Comp_5to3 c1_21(.X1(s0_0[21]), .X2(G[2][21-6]), .X3(G[3][21-9]), .X4(G[4][21-12]), .Ti(t1[20+1]),  .S(s1_0[21]), .C(c1_0[21+1]), .To(t1[21+1]));
    Comp_5to3 c1_22(.X1(s0_0[22]), .X2(c0_0[22]), .X3(G[2][22-6]), .X4(G[3][22-9]), .Ti(t1[21+1]),  .S(s1_0[22]), .C(c1_0[22+1]), .To(t1[22+1]));
    Comp_5to3 c1_23(.X1(s0_0[23]), .X2(c0_0[23]), .X3(G[2][23-6]), .X4(G[3][23-9]), .Ti(t1[22+1]),  .S(s1_0[23]), .C(c1_0[23+1]), .To(t1[23+1]));
    Comp_5to3 c1_24(.X1(s0_0[24]), .X2(c0_0[24]), .X3(G[3][24-9]), .X4(G[4][24-12]), .Ti(t1[23+1]),  .S(s1_0[24]), .C(c1_0[24+1]), .To(t1[24+1]));
    Comp_5to3 c1_25(.X1(s0_0[25]), .X2(c0_0[25]), .X3(G[3][25-9]), .X4(G[4][25-12]), .Ti(t1[24+1]),  .S(s1_0[25]), .C(c1_0[25+1]), .To(t1[25+1]));
    Comp_5to3 c1_26(.X1(s0_0[26]), .X2(c0_0[26]), .X3(G[3][26-9]), .X4(G[4][26-12]), .Ti(t1[25+1]),  .S(s1_0[26]), .C(c1_0[26+1]), .To(t1[26+1]));
    Comp_5to3 c1_27(.X1(s0_0[27]), .X2(c0_0[27]), .X3(G[3][27-9]), .X4(G[4][27-12]), .Ti(t1[26+1]),  .S(s1_0[27]), .C(c1_0[27+1]), .To(t1[27+1]));
    Comp_5to3 c1_28(.X1(s0_0[28]), .X2(c0_0[28]), .X3(G[3][28-9]), .X4(G[4][28-12]), .Ti(t1[27+1]),  .S(s1_0[28]), .C(c1_0[28+1]), .To(t1[28+1]));
    Comp_5to3 c1_29(.X1(s0_0[29]), .X2(c0_0[29]), .X3(G[3][29-9]), .X4(G[4][29-12]), .Ti(t1[28+1]),  .S(s1_0[29]), .C(c1_0[29+1]), .To(t1[29+1]));
    Comp_5to3 c1_30(.X1(s0_0[30]), .X2(c0_0[30]), .X3(G[3][30-9]), .X4(G[4][30-12]), .Ti(t1[29+1]),  .S(s1_0[30]), .C(c1_0[30+1]), .To(t1[30+1]));
    Comp_5to3 c1_31(.X1(s0_0[31]), .X2(c0_0[31]), .X3(G[3][31-9]), .X4(G[4][31-12]), .Ti(t1[30+1]),  .S(s1_0[31]), .C(c1_0[31+1]), .To(t1[31+1]));
    Comp_5to3 c1_32(.X1(~N[2]), .X2(c0_0[32]), .X3(G[3][32-9]), .X4(G[4][32-12]), .Ti(t1[31+1]),  .S(s1_0[32]), .C(c1_0[32+1]), .To(t1[32+1]));
    Comp_5to3 c1_33(.X1(1'b1), .X2(G[3][33-9]), .X3(G[4][33-12]), .X4(G[5][33-15]), .Ti(t1[32+1]),  .S(s1_0[33]), .C(c1_0[33+1]), .To(t1[33+1]));
    Comp_5to3 c1_34(.X1(1'b1), .X2(G[3][34-9]), .X3(G[4][34-12]), .X4(G[5][34-15]), .Ti(t1[33+1]),  .S(s1_0[34]), .C(c1_0[34+1]), .To(t1[34+1]));
    Comp_5to3 c1_35(.X1(~N[3]), .X2(G[4][35-12]), .X3(G[5][35-15]), .X4(G[6][35-18]), .Ti(t1[34+1]),  .S(s1_0[35]), .C(c1_0[35+1]), .To(t1[35+1]));
    Comp_4to2 c1_36(.X1(1'b1), .X2(G[4][36-12]), .X3(G[5][36-15]), .Ti(t1[35+1]),  .S(s1_0[36]), .C(c1_0[36+1]), .To(t1[36+1]));
    Comp_4to2 c1_37(.X1(1'b1), .X2(G[4][37-12]), .X3(G[5][37-15]), .Ti(t1[36+1]),  .S(s1_0[37]), .C(c1_0[37+1]), .To(t1[37+1]));
    FA c1_38(.A(~N[4]), .B(G[5][38-15]), .Ci(t1[37+1]),  .S(s1_0[38]), .Co(c1_0[38+1]));
    HA c1_39 (.A(1'b1), .B(G[5][39-15]), .S(s1_0[39]), .Co(c1_0[39+1]));
    HA c1_40 (.A(1'b1), .B(G[5][40-15]), .S(s1_0[40]), .Co(c1_0[40+1]));


	//******SECOND ROW OF COMPRESSORS IN THE SECOND LAYER******

    wire [34:18] s1_1;	//Sum outputs of the compressors (inputs of the next layer)
    wire [35:19] c1_1;	//Carry out of the compressors (inputs of the next layer)

    HA x1_18 (.A(G[4][18-12]), .B(G[5][18-15]), .S(s1_1[18]), .Co(c1_1[18+1]));
    HA x1_19 (.A(G[4][19-12]), .B(G[5][19-15]), .S(s1_1[19]), .Co(c1_1[19+1]));
    HA x1_20 (.A(G[4][20-12]), .B(G[5][20-15]), .S(s1_1[20]), .Co(c1_1[20+1]));
    FA x1_21 (.A(G[5][21-15]), .B(G[6][21-18]), .Ci(G[7][21-21]), .S(s1_1[21]), .Co(c1_1[21+1]));
    FA x1_22 (.A(G[4][22-12]), .B(G[5][22-15]), .Ci(G[6][22-18]), .S(s1_1[22]), .Co(c1_1[22+1]));
    FA x1_23 (.A(G[4][23-12]), .B(G[5][23-15]), .Ci(G[6][23-18]), .S(s1_1[23]), .Co(c1_1[23+1]));
    FA x1_24 (.A(G[5][24-15]), .B(G[6][24-18]), .Ci(G[7][24-21]), .S(s1_1[24]), .Co(c1_1[24+1]));
    FA x1_25 (.A(G[5][25-15]), .B(G[6][25-18]), .Ci(G[7][25-21]), .S(s1_1[25]), .Co(c1_1[25+1]));
    FA x1_26 (.A(G[5][26-15]), .B(G[6][26-18]), .Ci(G[7][26-21]), .S(s1_1[26]), .Co(c1_1[26+1]));
    FA x1_27 (.A(G[5][27-15]), .B(G[6][27-18]), .Ci(G[7][27-21]), .S(s1_1[27]), .Co(c1_1[27+1]));
    FA x1_28 (.A(G[5][28-15]), .B(G[6][28-18]), .Ci(G[7][28-21]), .S(s1_1[28]), .Co(c1_1[28+1]));
    FA x1_29 (.A(G[5][29-15]), .B(G[6][29-18]), .Ci(G[7][29-21]), .S(s1_1[29]), .Co(c1_1[29+1]));
    FA x1_30 (.A(G[5][30-15]), .B(G[6][30-18]), .Ci(G[7][30-21]), .S(s1_1[30]), .Co(c1_1[30+1]));
    FA x1_31 (.A(G[5][31-15]), .B(G[6][31-18]), .Ci(G[7][31-21]), .S(s1_1[31]), .Co(c1_1[31+1]));
    FA x1_32 (.A(G[5][32-15]), .B(G[6][32-18]), .Ci(G[7][32-21]), .S(s1_1[32]), .Co(c1_1[32+1]));
    HA x1_33 (.A(G[6][33-18]), .B(G[7][33-21]), .S(s1_1[33]), .Co(c1_1[33+1]));
    HA x1_34 (.A(G[6][34-18]), .B(G[7][34-21]), .S(s1_1[34]), .Co(c1_1[34+1]));


	//******THIRD LAYER******

    wire [46:6] s2_0;	//Sum outputs of the compressors (inputs of the next layer)
    wire [47:7] c2_0;	//Carry out of the compressors (inputs of the next layer)
    wire [44:10] t2;	//Intermediate T between compressors of te same layer

    HA c2_6 (.A(G[0][6]), .B(G[1][6-3]), .S(s2_0[6]), .Co(c2_0[6+1]));
    HA c2_7 (.A(G[0][7]), .B(G[1][7-3]), .S(s2_0[7]), .Co(c2_0[7+1]));
    HA c2_8 (.A(G[0][8]), .B(G[1][8-3]), .S(s2_0[8]), .Co(c2_0[8+1]));
    Comp_4to2 c2_9(.X1(G[0][9]), .X2(G[1][9-3]), .X3(G[2][9-6]), .Ti(G[3][9-9]),  .S(s2_0[9]), .C(c2_0[9+1]), .To(t2[9+1]));
    Comp_4to2 c2_10(.X1(G[0][10]), .X2(G[1][10-3]), .X3(G[2][10-6]), .Ti(t2[9+1]),  .S(s2_0[10]), .C(c2_0[10+1]), .To(t2[10+1]));
    Comp_4to2 c2_11(.X1(G[0][11]), .X2(G[1][11-3]), .X3(G[2][11-6]), .Ti(t2[10+1]),  .S(s2_0[11]), .C(c2_0[11+1]), .To(t2[11+1]));
    Comp_5to3 c2_12(.X1(s1_0[12]), .X2(G[2][12-6]), .X3(G[3][12-9]), .X4(G[4][12-12]), .Ti(t2[11+1]),  .S(s2_0[12]), .C(c2_0[12+1]), .To(t2[12+1]));
    Comp_5to3 c2_13(.X1(s1_0[13]), .X2(c1_0[13]), .X3(G[2][13-6]), .X4(G[3][13-9]), .Ti(t2[12+1]),  .S(s2_0[13]), .C(c2_0[13+1]), .To(t2[13+1]));
    Comp_5to3 c2_14(.X1(s1_0[14]), .X2(c1_0[14]), .X3(G[2][14-6]), .X4(G[3][14-9]), .Ti(t2[13+1]),  .S(s2_0[14]), .C(c2_0[14+1]), .To(t2[14+1]));
    Comp_5to3 c2_15(.X1(s1_0[15]), .X2(c1_0[15]), .X3(G[4][15-12]), .X4(G[5][15-15]), .Ti(t2[14+1]),  .S(s2_0[15]), .C(c2_0[15+1]), .To(t2[15+1]));
    Comp_5to3 c2_16(.X1(s1_0[16]), .X2(c1_0[16]), .X3(G[3][16-9]), .X4(G[4][16-12]), .Ti(t2[15+1]),  .S(s2_0[16]), .C(c2_0[16+1]), .To(t2[16+1]));
    Comp_5to3 c2_17(.X1(s1_0[17]), .X2(c1_0[17]), .X3(G[3][17-9]), .X4(G[4][17-12]), .Ti(t2[16+1]),  .S(s2_0[17]), .C(c2_0[17+1]), .To(t2[17+1]));
    Comp_5to3 c2_18(.X1(s1_0[18]), .X2(c1_0[18]), .X3(s1_1[18]), .X4(G[6][18-18]), .Ti(t2[17+1]),  .S(s2_0[18]), .C(c2_0[18+1]), .To(t2[18+1]));
    Comp_5to3 c2_19(.X1(s1_0[19]), .X2(c1_0[19]), .X3(s1_1[19]), .X4(c1_1[19]), .Ti(t2[18+1]),  .S(s2_0[19]), .C(c2_0[19+1]), .To(t2[19+1]));
    Comp_5to3 c2_20(.X1(s1_0[20]), .X2(c1_0[20]), .X3(s1_1[20]), .X4(c1_1[20]), .Ti(t2[19+1]),  .S(s2_0[20]), .C(c2_0[20+1]), .To(t2[20+1]));
    Comp_5to3 c2_21(.X1(s1_0[21]), .X2(c1_0[21]), .X3(s1_1[21]), .X4(c1_1[21]), .Ti(t2[20+1]),  .S(s2_0[21]), .C(c2_0[21+1]), .To(t2[21+1]));
    Comp_5to3 c2_22(.X1(s1_0[22]), .X2(c1_0[22]), .X3(s1_1[22]), .X4(c1_1[22]), .Ti(t2[21+1]),  .S(s2_0[22]), .C(c2_0[22+1]), .To(t2[22+1]));
    Comp_5to3 c2_23(.X1(s1_0[23]), .X2(c1_0[23]), .X3(s1_1[23]), .X4(c1_1[23]), .Ti(t2[22+1]),  .S(s2_0[23]), .C(c2_0[23+1]), .To(t2[23+1]));
    Comp_5to3 c2_24(.X1(s1_0[24]), .X2(c1_0[24]), .X3(s1_1[24]), .X4(c1_1[24]), .Ti(t2[23+1]),  .S(s2_0[24]), .C(c2_0[24+1]), .To(t2[24+1]));
    Comp_5to3 c2_25(.X1(s1_0[25]), .X2(c1_0[25]), .X3(s1_1[25]), .X4(c1_1[25]), .Ti(t2[24+1]),  .S(s2_0[25]), .C(c2_0[25+1]), .To(t2[25+1]));
    Comp_5to3 c2_26(.X1(s1_0[26]), .X2(c1_0[26]), .X3(s1_1[26]), .X4(c1_1[26]), .Ti(t2[25+1]),  .S(s2_0[26]), .C(c2_0[26+1]), .To(t2[26+1]));
    Comp_5to3 c2_27(.X1(s1_0[27]), .X2(c1_0[27]), .X3(s1_1[27]), .X4(c1_1[27]), .Ti(t2[26+1]),  .S(s2_0[27]), .C(c2_0[27+1]), .To(t2[27+1]));
    Comp_5to3 c2_28(.X1(s1_0[28]), .X2(c1_0[28]), .X3(s1_1[28]), .X4(c1_1[28]), .Ti(t2[27+1]),  .S(s2_0[28]), .C(c2_0[28+1]), .To(t2[28+1]));
    Comp_5to3 c2_29(.X1(s1_0[29]), .X2(c1_0[29]), .X3(s1_1[29]), .X4(c1_1[29]), .Ti(t2[28+1]),  .S(s2_0[29]), .C(c2_0[29+1]), .To(t2[29+1]));
    Comp_5to3 c2_30(.X1(s1_0[30]), .X2(c1_0[30]), .X3(s1_1[30]), .X4(c1_1[30]), .Ti(t2[29+1]),  .S(s2_0[30]), .C(c2_0[30+1]), .To(t2[30+1]));
    Comp_5to3 c2_31(.X1(s1_0[31]), .X2(c1_0[31]), .X3(s1_1[31]), .X4(c1_1[31]), .Ti(t2[30+1]),  .S(s2_0[31]), .C(c2_0[31+1]), .To(t2[31+1]));
    Comp_5to3 c2_32(.X1(s1_0[32]), .X2(c1_0[32]), .X3(s1_1[32]), .X4(c1_1[32]), .Ti(t2[31+1]),  .S(s2_0[32]), .C(c2_0[32+1]), .To(t2[32+1]));
    Comp_5to3 c2_33(.X1(s1_0[33]), .X2(c1_0[33]), .X3(s1_1[33]), .X4(c1_1[33]), .Ti(t2[32+1]),  .S(s2_0[33]), .C(c2_0[33+1]), .To(t2[33+1]));
    Comp_5to3 c2_34(.X1(s1_0[34]), .X2(c1_0[34]), .X3(s1_1[34]), .X4(c1_1[34]), .Ti(t2[33+1]),  .S(s2_0[34]), .C(c2_0[34+1]), .To(t2[34+1]));
    Comp_5to3 c2_35(.X1(s1_0[35]), .X2(c1_0[35]), .X3(G[7][35-21]), .X4(c1_1[35]), .Ti(t2[34+1]),  .S(s2_0[35]), .C(c2_0[35+1]), .To(t2[35+1]));
    Comp_5to3 c2_36(.X1(s1_0[36]), .X2(c1_0[36]), .X3(G[6][36-18]), .X4(G[7][36-21]), .Ti(t2[35+1]),  .S(s2_0[36]), .C(c2_0[36+1]), .To(t2[36+1]));
    Comp_5to3 c2_37(.X1(s1_0[37]), .X2(c1_0[37]), .X3(G[6][37-18]), .X4(G[7][37-21]), .Ti(t2[36+1]),  .S(s2_0[37]), .C(c2_0[37+1]), .To(t2[37+1]));
    Comp_5to3 c2_38(.X1(s1_0[38]), .X2(c1_0[38]), .X3(G[6][38-18]), .X4(G[7][38-21]), .Ti(t2[37+1]),  .S(s2_0[38]), .C(c2_0[38+1]), .To(t2[38+1]));
    Comp_5to3 c2_39(.X1(s1_0[39]), .X2(c1_0[39]), .X3(G[6][39-18]), .X4(G[7][39-21]), .Ti(t2[38+1]),  .S(s2_0[39]), .C(c2_0[39+1]), .To(t2[39+1]));
    Comp_5to3 c2_40(.X1(s1_0[40]), .X2(c1_0[40]), .X3(G[6][40-18]), .X4(G[7][40-21]), .Ti(t2[39+1]),  .S(s2_0[40]), .C(c2_0[40+1]), .To(t2[40+1]));
    Comp_5to3 c2_41(.X1(~N[5]), .X2(c1_0[41]), .X3(G[6][41-18]), .X4(G[7][41-21]), .Ti(t2[40+1]),  .S(s2_0[41]), .C(c2_0[41+1]), .To(t2[41+1]));
    Comp_4to2 c2_42(.X1(1'b1), .X2(G[6][42-18]), .X3(G[7][42-21]), .Ti(t2[41+1]),  .S(s2_0[42]), .C(c2_0[42+1]), .To(t2[42+1]));
    Comp_4to2 c2_43(.X1(1'b1), .X2(G[6][43-18]), .X3(G[7][43-21]), .Ti(t2[42+1]),  .S(s2_0[43]), .C(c2_0[43+1]), .To(t2[43+1]));
    FA c2_44 (.A(~N[6]), .B(G[7][44-21]), .Ci(t2[43+1]), .S(s2_0[44]), .Co(c2_0[44+1]));
    HA c2_45 (.A(1'b1), .B(G[7][45-21]), .S(s2_0[45]), .Co(c2_0[45+1]));
    HA c2_46 (.A(1'b1), .B(G[7][46-21]), .S(s2_0[46]), .Co(c2_0[46+1]));


	//******FOURTH LAYER******

    wire [49:3] s3_0;	//Sum outputs of the compressors (inputs of the next layer)
    wire [50:4] c3_0;	//Carry out of the compressors (inputs of the next layer)
    
    HA c3_3 (.A(G[0][3]), .B(G[1][3-3]), .S(s3_0[3]), .Co(c3_0[3+1]));
    HA c3_4 (.A(G[0][4]), .B(G[1][4-3]), .S(s3_0[4]), .Co(c3_0[4+1]));
    HA c3_5 (.A(G[0][5]), .B(G[1][5-3]), .S(s3_0[5]), .Co(c3_0[5+1]));
    FA c3_6 (.A(s2_0[6]), .B(G[2][6-6]), .Ci(N[2]), .S(s3_0[6]), .Co(c3_0[6+1]));
    FA c3_7 (.A(s2_0[7]), .B(c2_0[7]), .Ci(G[2][7-6]), .S(s3_0[7]), .Co(c3_0[7+1]));
    FA c3_8 (.A(s2_0[8]), .B(c2_0[8]), .Ci(G[2][8-6]), .S(s3_0[8]), .Co(c3_0[8+1]));
    FA c3_9 (.A(s2_0[9]), .B(c2_0[9]), .Ci(N[3]), .S(s3_0[9]), .Co(c3_0[9+1]));
    FA c3_10 (.A(s2_0[10]), .B(c2_0[10]), .Ci(G[3][10-9]), .S(s3_0[10]), .Co(c3_0[10+1]));
    FA c3_11 (.A(s2_0[11]), .B(c2_0[11]), .Ci(G[3][11-9]), .S(s3_0[11]), .Co(c3_0[11+1]));
    FA c3_12 (.A(s2_0[12]), .B(c2_0[12]), .Ci(N[4]), .S(s3_0[12]), .Co(c3_0[12+1]));
    FA c3_13 (.A(s2_0[13]), .B(c2_0[13]), .Ci(G[4][13-12]), .S(s3_0[13]), .Co(c3_0[13+1]));
    FA c3_14 (.A(s2_0[14]), .B(c2_0[14]), .Ci(G[4][14-12]), .S(s3_0[14]), .Co(c3_0[14+1]));
    FA c3_15 (.A(s2_0[15]), .B(c2_0[15]), .Ci(N[5]), .S(s3_0[15]), .Co(c3_0[15+1]));
    FA c3_16 (.A(s2_0[16]), .B(c2_0[16]), .Ci(G[5][16-15]), .S(s3_0[16]), .Co(c3_0[16+1]));
    FA c3_17 (.A(s2_0[17]), .B(c2_0[17]), .Ci(G[5][17-15]), .S(s3_0[17]), .Co(c3_0[17+1]));
    FA c3_18 (.A(s2_0[18]), .B(c2_0[18]), .Ci(N[6]), .S(s3_0[18]), .Co(c3_0[18+1]));
    FA c3_19 (.A(s2_0[19]), .B(c2_0[19]), .Ci(G[6][19-18]), .S(s3_0[19]), .Co(c3_0[19+1]));
    FA c3_20 (.A(s2_0[20]), .B(c2_0[20]), .Ci(G[6][20-18]), .S(s3_0[20]), .Co(c3_0[20+1]));
    FA c3_21 (.A(s2_0[21]), .B(c2_0[21]), .Ci(N[7]), .S(s3_0[21]), .Co(c3_0[21+1]));
    FA c3_22 (.A(s2_0[22]), .B(c2_0[22]), .Ci(G[7][22-21]), .S(s3_0[22]), .Co(c3_0[22+1]));
    FA c3_23 (.A(s2_0[23]), .B(c2_0[23]), .Ci(G[7][23-21]), .S(s3_0[23]), .Co(c3_0[23+1]));
    FA c3_24 (.A(s2_0[24]), .B(c2_0[24]), .Ci(G[8][24-24]), .S(s3_0[24]), .Co(c3_0[24+1]));
    FA c3_25 (.A(s2_0[25]), .B(c2_0[25]), .Ci(G[8][25-24]), .S(s3_0[25]), .Co(c3_0[25+1]));
    FA c3_26 (.A(s2_0[26]), .B(c2_0[26]), .Ci(G[8][26-24]), .S(s3_0[26]), .Co(c3_0[26+1]));
    FA c3_27 (.A(s2_0[27]), .B(c2_0[27]), .Ci(G[8][27-24]), .S(s3_0[27]), .Co(c3_0[27+1]));
    FA c3_28 (.A(s2_0[28]), .B(c2_0[28]), .Ci(G[8][28-24]), .S(s3_0[28]), .Co(c3_0[28+1]));
    FA c3_29 (.A(s2_0[29]), .B(c2_0[29]), .Ci(G[8][29-24]), .S(s3_0[29]), .Co(c3_0[29+1]));
    FA c3_30 (.A(s2_0[30]), .B(c2_0[30]), .Ci(G[8][30-24]), .S(s3_0[30]), .Co(c3_0[30+1]));
    FA c3_31 (.A(s2_0[31]), .B(c2_0[31]), .Ci(G[8][31-24]), .S(s3_0[31]), .Co(c3_0[31+1]));
    FA c3_32 (.A(s2_0[32]), .B(c2_0[32]), .Ci(G[8][32-24]), .S(s3_0[32]), .Co(c3_0[32+1]));
    FA c3_33 (.A(s2_0[33]), .B(c2_0[33]), .Ci(G[8][33-24]), .S(s3_0[33]), .Co(c3_0[33+1]));
    FA c3_34 (.A(s2_0[34]), .B(c2_0[34]), .Ci(G[8][34-24]), .S(s3_0[34]), .Co(c3_0[34+1]));
    FA c3_35 (.A(s2_0[35]), .B(c2_0[35]), .Ci(G[8][35-24]), .S(s3_0[35]), .Co(c3_0[35+1]));
    FA c3_36 (.A(s2_0[36]), .B(c2_0[36]), .Ci(G[8][36-24]), .S(s3_0[36]), .Co(c3_0[36+1]));
    FA c3_37 (.A(s2_0[37]), .B(c2_0[37]), .Ci(G[8][37-24]), .S(s3_0[37]), .Co(c3_0[37+1]));
    FA c3_38 (.A(s2_0[38]), .B(c2_0[38]), .Ci(G[8][38-24]), .S(s3_0[38]), .Co(c3_0[38+1]));
    FA c3_39 (.A(s2_0[39]), .B(c2_0[39]), .Ci(G[8][39-24]), .S(s3_0[39]), .Co(c3_0[39+1]));
    FA c3_40 (.A(s2_0[40]), .B(c2_0[40]), .Ci(G[8][40-24]), .S(s3_0[40]), .Co(c3_0[40+1]));
    FA c3_41 (.A(s2_0[41]), .B(c2_0[41]), .Ci(G[8][41-24]), .S(s3_0[41]), .Co(c3_0[41+1]));
    FA c3_42 (.A(s2_0[42]), .B(c2_0[42]), .Ci(G[8][42-24]), .S(s3_0[42]), .Co(c3_0[42+1]));
    FA c3_43 (.A(s2_0[43]), .B(c2_0[43]), .Ci(G[8][43-24]), .S(s3_0[43]), .Co(c3_0[43+1]));
    FA c3_44 (.A(s2_0[44]), .B(c2_0[44]), .Ci(G[8][44-24]), .S(s3_0[44]), .Co(c3_0[44+1]));
    FA c3_45 (.A(s2_0[45]), .B(c2_0[45]), .Ci(G[8][45-24]), .S(s3_0[45]), .Co(c3_0[45+1]));
    FA c3_46 (.A(s2_0[46]), .B(c2_0[46]), .Ci(G[8][46-24]), .S(s3_0[46]), .Co(c3_0[46+1]));
    FA c3_47 (.A(~N[7]), .B(c2_0[47]), .Ci(G[8][47-24]), .S(s3_0[47]), .Co(c3_0[47+1]));
    HA c3_48 (.A(1'b1), .B(G[8][48-24]), .S(s3_0[48]), .Co(c3_0[48+1]));
    HA c3_49 (.A(1'b1), .B(G[8][49-24]), .S(s3_0[49]), .Co(c3_0[49+1]));

    
    //******SUM OF THE FINAL TWO OPERANDS******

    wire [47:0] A;	//First operand
    wire [47:0] B;	//Second operand

    assign A = {s3_0[47:3], G[0][2:0]};
    assign B = {c3_0[47:4], N[1], 2'b0, N[0]};
    assign Z = A + B;	//Final addition
   
endmodule
